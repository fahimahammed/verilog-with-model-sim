module xnor_gate(A, B, Y);
input A, B;
output Y;

xnor(Y, A, B);


endmodule
