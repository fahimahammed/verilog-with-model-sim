module or_gate(A, B, Y);
input A, B;
output Y;
assign Y = A || B;
endmodule
